`timescale 1ns/1ps

`include "../rtl/_parameter.v"

// g = n + 1, lambda * mu = 1 (mod n)

module paillier_demo_overall_top_tb();
    reg clk;
    reg rst_n;
    parameter [15:0] width  = 4096;
    reg [(width - 1):0] c, c1, c2, m, r, n, exp_n, g, mu, lambda;
    reg [3:0] state;
    reg  go;
    wire done;
    wire [(width - 1):0] result;

    initial begin
        
        $dumpfile("rsa4k.vcd");
  		$dumpvars(0);

        clk = 0;

        #10
        rst_n = 0;
        #10
        rst_n = 1;
        go = 0;
        state = 4'b0000;

       
        $display("Test Case begin: 1. encry ");
        m = 4096'd914850650102228807940294227641046146757155842252766216264036753726262461423906917348160457992600443343560250435223363421123229695023423749360952614842508876914842205991852825524617900409935435880783844922223497593605542245610386263846464261837145187897364026566090205971196227826138905573642115708886515076561984749472544338169455942906187552477104159453455785061156306462028550638591670446353085326639557811752581457786411393004696664147460330131698788674030107577879239046357400994355357847699891799743490606164589910112977127754536023351516070966196151585029312678131220203158479344495472793961393548277830957646;
        r = 4096'd13407807929942597099574024998205846127479365820592393377723561443721764030073546976801874298166903427690031858186486050853753882811946569946433649006084096;
        n = 4096'd105246209408553047249848144100971688447826338579860315035513589711994872594953240247665410233278147844418006191557867876488977231998217690408511034339655074295010618073191295602931120109906709329940570153998669271048141423037028763471597408964025339740750277073920283582024037723473789898757244183003510744273;
        exp_n = 4096'd11076764594868999963804378401762617032843845914649700042044765379608002766441553535933585621427077945799258757592198128515613386910620126399332596165349860671405120483761974197000953867034096281236352265483748686430214197439487252724102734880261418131327993299372132238825571350317786056455641474066335045244448512169618316475851288926428399204545257762385330789010317773882105633978526358747499887965702270923938320697026162103401726008956494892259602926066905782698197629045020010449581733096982320383567668720148264679453234866970737732228497009815739838198190906481283943394788551792671978665471953243350402298529;
        g = 4096'd8383956268357347042308682846077637595761898737863014975857279871963667677465447427985078675253088055444944571431239397408949190232821295137186212970282539898877422547596549894449412046907720369833916647961752948691784986793149190411225628099315102358423890701615033737070008694741863927638590386230140631266390777896485325549852289518453249186221364520016733929948352748329599727651400038064727189420654239799168757040159078778674164200827938559528814224461442698159297561704067050344546980355352878912876018089595800835871442015272875580704492908052915012670604635358889243148195301570773332980543961426680671212102;

        state = 4'b0001;

        go = 1;
        #10
        wait(done);
        $display("[paillier_demo_overall_top_tb.v]result: \n0x%x",result);
        wait(!done);
        go = 0;
        
        #5
        #10
        rst_n = 0;
        #10
        rst_n = 1;
        
        
        $display("Test Case begin: 2. decry ");    
        c = 4096'd33524;
        lambda = 4096'd90;
        n = 4096'd209;
        exp_n = 4096'd43681;
        mu = 4096'd72;

        state = 4'b0010;

        go = 1;
        #10
        wait(done);
        $display("[paillier_demo_top_tb.v]result: \n0x%x",result);    
        wait(!done);

        go = 0;
        
        #10
        rst_n = 0;
        #10
        rst_n = 1;

        
        $display("Test Case begin: 3. homo add ");
        c1 = 4096'd226;
        c2 = 4096'd3409;
        n = 4096'd209;
        exp_n = 4096'd43681;

        state = 4'b0100;
        
        go = 1;
        #10
        wait(done);
        $display("[paillier_demo_overall_top_tb.v]result: \n0x%x",result);
        wait(!done);
        
        go = 0;
        
        #10
        rst_n = 0;
        #10
        rst_n = 1;

        
        $display("Test Case begin: 4. homo mul ");
        c = 4096'd226;
        m = 4096'd10;
        n = 4096'd209;
        exp_n = 4096'd43681;


        state = 4'b1000;

        go = 1;
        #10
        wait(done);
        $display("[paillier_demo_overall_top_tb.v]result: \n0x%x",result);
        wait(!done);
        
        $finish;

    end


    always begin
        #5 clk = ~clk;
    end

    paillier_demo_overall_top#(
        .RSA_WIDTH(4096),
        .DATA_WIDTH(128),
        .DATA_NUMBER(32)
    ) 
    paillier_demo_overall_top_u(
        .clk(clk),
        .rst_n(rst_n),
        .go(go),
        .m(m),
        .r(r),
        .c(c),
        .c1(c1),
        .c2(c2),
        .n(n),
        .exp_n(exp_n),
        .g(g),
        .lambda(lambda),
        .mu(mu),
        .state(state),
        .result(result),
        .done(done)
    );

endmodule